
ioadsjkj`
