i am naveen
getting started to github
