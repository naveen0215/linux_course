i am naveen
getting started to github
module tb;
logic a,b;
logic out;
assign out = a&b;
endmodule
