module tb;
inputs a,b;
output sum;
assign sum = a+b;
endmodule

