module vinay;

endmoduele
