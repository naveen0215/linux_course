I AM NAVEEN
NOW TO LEARN THE GITHUB COMMANDS
