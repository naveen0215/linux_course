nsjdnscnaskn
